`timescale 1ns / 1ps

// general purpose FIFO module

module FIFO #(parameter
  // TODO
) (
  // TODO
);

  // TODO

endmodule // FIFO
