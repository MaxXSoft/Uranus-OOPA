`timescale 1ns / 1ps

module Core(
  input clk,
  input rst,
  input [4:0] intr
);

//

endmodule // Core
